library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Gray_Counter_Tb is 
end entity;

architecture sim of Gray_Counter_Tb is 

-- Operational signals 
signal rst : std_logic := '0';
signal eneable : std_logic := '0';
signal clk	: std_logic := '0';
signal some_signal : std_logic := '0';

-- Constans
Constant Ctr_Size 	: natural := 8;
constant clk_period : time := 1 ns;


signal Nx 	: std_logic_vector(Ctr_Size - 1 downto 0);

procedure Wait_Raising_Edges (signal clk : in std_logic; n : integer) is 
begin
	for i in 1 to n loop
		wait until rising_edge(clk);
	end loop;

end procedure;

begin	
	rst <= '1', '0' after 2 ns;
	eneable <= '0', '1' after 1 ns;

	-- Instance device under test
	DUT: entity work.Gray_Counter(rtl)
	generic map(
	 WIDTH => Ctr_Size 
	)
	port map(
		clk	=>	clk,
	        reset	=>	rst,
	 	eneable	=>	eneable,
	       	gray_count =>	Nx
	);
	
	clk_process :process
   	begin
    		clk <= '0';
    		wait for clk_period/2; 
    		clk <= '1';
    		wait for clk_period/2;
   	end process;

	--some_stim_proc : process begin
	--	some_signal <= '0';
	-- 	Wait_Raising_Edges(clk,900);
	--	some_signal <= '1';
	-- 	Wait_Raising_Edges(clk,100);
	--	wait;	
	--end process;

end architecture;


 
